`timescale 1ns / 10ps

module SubBytes(matrix_in, matrix_out);
input wire [7:0] matrix_in;     // 8-bit input vector
output wire [7:0] matrix_out;   // 8-bit output vector

// Declare 16x16 array of 8bit 
reg [7:0] lookupTable [0:15][0:15];

// Manual SBOX Lookup Table
initial begin
    lookupTable[0][0] <= 8'h63; lookupTable[0][1] <= 8'h7c; lookupTable[0][2] = 8'h77; lookupTable[0][3] <= 8'h7b; lookupTable[0][4] <= 8'hf2; lookupTable[0][5] <= 8'h6b; lookupTable[0][6] = 8'h6f; lookupTable[0][7] <= 8'hc5; lookupTable[0][8] <= 8'h30; lookupTable[0][9] <= 8'h01; lookupTable[0][10] <= 8'h67; lookupTable[0][11] = 8'h2b; lookupTable[0][12] <= 8'hfe; lookupTable[0][13] <= 8'hd7; lookupTable[0][14] <= 8'hab; lookupTable[0][15] <= 8'h76; 
    lookupTable[1][0] <= 8'hca; lookupTable[1][1] <= 8'h82; lookupTable[1][2] = 8'hc9; lookupTable[1][3] <= 8'h7d; lookupTable[1][4] <= 8'hfa; lookupTable[1][5] <= 8'h59; lookupTable[1][6] = 8'h47; lookupTable[1][7] <= 8'hf0; lookupTable[1][8] <= 8'had; lookupTable[1][9] <= 8'hd4; lookupTable[1][10] <= 8'ha2; lookupTable[1][11] = 8'haf; lookupTable[1][12] <= 8'h9c; lookupTable[1][13] <= 8'ha4; lookupTable[1][14] <= 8'h72; lookupTable[1][15] <= 8'hc0; 
    lookupTable[2][0] <= 8'hb7; lookupTable[2][1] <= 8'hfd; lookupTable[2][2] = 8'h93; lookupTable[2][3] <= 8'h26; lookupTable[2][4] <= 8'h36; lookupTable[2][5] <= 8'h3f; lookupTable[2][6] = 8'hf7; lookupTable[2][7] <= 8'hcc; lookupTable[2][8] <= 8'h34; lookupTable[2][9] <= 8'ha5; lookupTable[2][10] <= 8'he5; lookupTable[2][11] = 8'hf1; lookupTable[2][12] <= 8'h71; lookupTable[2][13] <= 8'hd8; lookupTable[2][14] <= 8'h31; lookupTable[2][15] <= 8'h15; 
    lookupTable[3][0] <= 8'h04; lookupTable[3][1] <= 8'hc7; lookupTable[3][2] = 8'h23; lookupTable[3][3] <= 8'hc3; lookupTable[3][4] <= 8'h18; lookupTable[3][5] <= 8'h96; lookupTable[3][6] = 8'h05; lookupTable[3][7] <= 8'h9a; lookupTable[3][8] <= 8'h07; lookupTable[3][9] <= 8'h12; lookupTable[3][10] <= 8'h80; lookupTable[3][11] = 8'he2; lookupTable[3][12] <= 8'heb; lookupTable[3][13] <= 8'h27; lookupTable[3][14] <= 8'hb2; lookupTable[3][15] <= 8'h75; 
    lookupTable[4][0] <= 8'h09; lookupTable[4][1] <= 8'h83; lookupTable[4][2] = 8'h2c; lookupTable[4][3] <= 8'h1a; lookupTable[4][4] <= 8'h1b; lookupTable[4][5] <= 8'h6e; lookupTable[4][6] = 8'h5a; lookupTable[4][7] <= 8'ha0; lookupTable[4][8] <= 8'h52; lookupTable[4][9] <= 8'h3b; lookupTable[4][10] <= 8'hd6; lookupTable[4][11] = 8'hb3; lookupTable[4][12] <= 8'h29; lookupTable[4][13] <= 8'he3; lookupTable[4][14] <= 8'h2f; lookupTable[4][15] <= 8'h84;
    lookupTable[5][0] <= 8'h53; lookupTable[5][1] <= 8'hd1; lookupTable[5][2] = 8'h00; lookupTable[5][3] <= 8'hed; lookupTable[5][4] <= 8'h20; lookupTable[5][5] <= 8'hfc; lookupTable[5][6] = 8'hb1; lookupTable[5][7] <= 8'h5b; lookupTable[5][8] <= 8'h6a; lookupTable[5][9] <= 8'hcb; lookupTable[5][10] <= 8'hbe; lookupTable[5][11] = 8'h39; lookupTable[5][12] <= 8'h4a; lookupTable[5][13] <= 8'h4c; lookupTable[5][14] <= 8'h58; lookupTable[5][15] <= 8'hcf;
    lookupTable[6][0] <= 8'hd0; lookupTable[6][1] <= 8'hef; lookupTable[6][2] = 8'haa; lookupTable[6][3] <= 8'hfb; lookupTable[6][4] <= 8'h43; lookupTable[6][5] <= 8'h4d; lookupTable[6][6] = 8'h33; lookupTable[6][7] <= 8'h85; lookupTable[6][8] <= 8'h45; lookupTable[6][9] <= 8'hf9; lookupTable[6][10] <= 8'h02; lookupTable[6][11] = 8'h7f; lookupTable[6][12] <= 8'h50; lookupTable[6][13] <= 8'h3c; lookupTable[6][14] <= 8'h9f; lookupTable[6][15] <= 8'ha8;
    lookupTable[7][0] <= 8'h51; lookupTable[7][1] <= 8'ha3; lookupTable[7][2] = 8'h40; lookupTable[7][3] <= 8'h8f; lookupTable[7][4] <= 8'h92; lookupTable[7][5] <= 8'h9d; lookupTable[7][6] = 8'h38; lookupTable[7][7] <= 8'hf5; lookupTable[7][8] <= 8'hbc; lookupTable[7][9] <= 8'hb6; lookupTable[7][10] <= 8'hda; lookupTable[7][11] = 8'h21; lookupTable[7][12] <= 8'h10; lookupTable[7][13] <= 8'hff; lookupTable[7][14] <= 8'hf3; lookupTable[7][15] <= 8'hd2;
    lookupTable[8][0] <= 8'hcd; lookupTable[8][1] <= 8'h0c; lookupTable[8][2] = 8'h13; lookupTable[8][3] <= 8'hec; lookupTable[8][4] <= 8'h5f; lookupTable[8][5] <= 8'h97; lookupTable[8][6] = 8'h44; lookupTable[8][7] <= 8'h17; lookupTable[8][8] <= 8'hc4; lookupTable[8][9] <= 8'ha7; lookupTable[8][10] <= 8'h7e; lookupTable[8][11] = 8'h3d; lookupTable[8][12] <= 8'h64; lookupTable[8][13] <= 8'h5d; lookupTable[8][14] <= 8'h19; lookupTable[8][15] <= 8'h73;
    lookupTable[9][0] <= 8'h60; lookupTable[9][1] <= 8'h81; lookupTable[9][2] = 8'h4f; lookupTable[9][3] <= 8'hdc; lookupTable[9][4] <= 8'h22; lookupTable[9][5] <= 8'h2a; lookupTable[9][6] = 8'h90; lookupTable[9][7] <= 8'h88; lookupTable[9][8] <= 8'h46; lookupTable[9][9] <= 8'hee; lookupTable[9][10] <= 8'hb8; lookupTable[9][11] = 8'h14; lookupTable[9][12] <= 8'hde; lookupTable[9][13] <= 8'h5e; lookupTable[9][14] <= 8'h0b; lookupTable[9][15] <= 8'hdb;
    lookupTable[10][0] <= 8'he0; lookupTable[10][1] <= 8'h32; lookupTable[10][2] = 8'h3a; lookupTable[10][3] <= 8'h0a; lookupTable[10][4] <= 8'h49; lookupTable[10][5] <= 8'h06; lookupTable[10][6] = 8'h24; lookupTable[10][7] <= 8'h5c; lookupTable[10][8] <= 8'hc2; lookupTable[10][9] <= 8'hd3; lookupTable[10][10] = 8'hac; lookupTable[10][11] <= 8'h62; lookupTable[10][12] <= 8'h91; lookupTable[10][13] <= 8'h95; lookupTable[10][14] <= 8'he4; lookupTable[10][15] <= 8'h79;
    lookupTable[11][0] <= 8'he7; lookupTable[11][1] <= 8'hc8; lookupTable[11][2] = 8'h37; lookupTable[11][3] <= 8'h6d; lookupTable[11][4] <= 8'h8d; lookupTable[11][5] <= 8'hd5; lookupTable[11][6] = 8'h4e; lookupTable[11][7] <= 8'ha9; lookupTable[11][8] <= 8'h6c; lookupTable[11][9] <= 8'h56; lookupTable[11][10] = 8'hf4; lookupTable[11][11] <= 8'hea; lookupTable[11][12] <= 8'h65; lookupTable[11][13] <= 8'h7a; lookupTable[11][14] <= 8'hae; lookupTable[11][15] <= 8'h08;
    lookupTable[12][0] <= 8'hba; lookupTable[12][1] <= 8'h78; lookupTable[12][2] = 8'h25; lookupTable[12][3] <= 8'h2e; lookupTable[12][4] <= 8'h1c; lookupTable[12][5] <= 8'ha6; lookupTable[12][6] = 8'hb4; lookupTable[12][7] <= 8'hc6; lookupTable[12][8] <= 8'he8; lookupTable[12][9] <= 8'hdd; lookupTable[12][10] = 8'h74; lookupTable[12][11] <= 8'h1f; lookupTable[12][12] <= 8'h4b; lookupTable[12][13] <= 8'hbd; lookupTable[12][14] <= 8'h8b; lookupTable[12][15] <= 8'h8a;
    lookupTable[13][0] <= 8'h70; lookupTable[13][1] <= 8'h3e; lookupTable[13][2] = 8'hb5; lookupTable[13][3] <= 8'h66; lookupTable[13][4] <= 8'h48; lookupTable[13][5] <= 8'h03; lookupTable[13][6] = 8'hf6; lookupTable[13][7] <= 8'h0e; lookupTable[13][8] <= 8'h61; lookupTable[13][9] <= 8'h35; lookupTable[13][10] = 8'h57; lookupTable[13][11] <= 8'hb9; lookupTable[13][12] <= 8'h86; lookupTable[13][13] <= 8'hc1; lookupTable[13][14] <= 8'h1d; lookupTable[13][15] <= 8'h9e;
    lookupTable[14][0] <= 8'he1; lookupTable[14][1] <= 8'hf8; lookupTable[14][2] = 8'h98; lookupTable[14][3] <= 8'h11; lookupTable[14][4] <= 8'h69; lookupTable[14][5] <= 8'hd9; lookupTable[14][6] = 8'h8e; lookupTable[14][7] <= 8'h94; lookupTable[14][8] <= 8'h9b; lookupTable[14][9] <= 8'h1e; lookupTable[14][10] = 8'h87; lookupTable[14][11] <= 8'he9; lookupTable[14][12] <= 8'hce; lookupTable[14][13] <= 8'h55; lookupTable[14][14] <= 8'h28; lookupTable[14][15] <= 8'hdf;
    lookupTable[15][0] <= 8'h8c; lookupTable[15][1] <= 8'ha1; lookupTable[15][2] = 8'h89; lookupTable[15][3] <= 8'h0d; lookupTable[15][4] <= 8'hbf; lookupTable[15][5] <= 8'he6; lookupTable[15][6] = 8'h42; lookupTable[15][7] <= 8'h68; lookupTable[15][8] <= 8'h41; lookupTable[15][9] <= 8'h99; lookupTable[15][10] = 8'h2d; lookupTable[15][11] <= 8'h0f; lookupTable[15][12] <= 8'hb0; lookupTable[15][13] <= 8'h54; lookupTable[15][14] <= 8'hbb; lookupTable[15][15] <= 8'h16;
end

assign matrix_out = lookupTable[matrix_in[7:4]][matrix_in[3:0]];
endmodule